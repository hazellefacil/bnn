library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity bnn is
  port(
  
		);
end bnn;

-- Architecture part of the description

architecture behavioural of bnn is


begin
	
end behavioural;