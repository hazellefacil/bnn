library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity binMatxbinVec is
  port(
  
		);
end binMatxbinVec;

-- Architecture part of the description

architecture behavioural of binMatxbinVec is


begin
	
end behavioural;