library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity popcnt is
  port(
  
		);
end popcnt;

-- Architecture part of the description

architecture behavioural of popcnt is


begin
	
end behavioural;