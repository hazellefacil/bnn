library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity full_adder is
  port(
  
		);
end full_adder;

-- Architecture part of the description

architecture behavioural of full_adder is


begin
	
end behavioural;