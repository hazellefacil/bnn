library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity binMatxfullPrecisionVec is
  port(
  
		);
end binMatxfullPrecisionVec;

-- Architecture part of the description

architecture behavioural of binMatxfullPrecisionVec is


begin
	
end behavioural;