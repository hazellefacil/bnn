library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity x_norm is
  port(
  
		);
end x_norm;

-- Architecture part of the description

architecture behavioural of x_norm is


begin
	
end behavioural;