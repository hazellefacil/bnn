library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity Bn is
  port(
  
		);
end Bn;

-- Architecture part of the description

architecture behavioural of Bn is


begin
	
end behavioural;