LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY popcnt_128 IS
	GENERIC(N	: NATURAL := 128); 
	PORT(INPUT 	: IN  STD_LOGIC_VECTOR(N-1 downto 0);
		SUM		: OUT INTEGER := 0;
		DONE		: OUT STD_LOGIC := '0'); 
END popcnt_128;

ARCHITECTURE RTL OF popcnt_128 IS	 
	
BEGIN	

	PROCESS(INPUT) 
		VARIABLE tempSUM	:	INTEGER := 0;
		CONSTANT ZERO		:	INTEGER := 0;
		CONSTANT COUNT_MAX	:	INTEGER := N - 1;
	BEGIN 

		DONE <= '0';
		tempSUM := 0;
		
		FOR COUNT IN 0 TO COUNT_MAX LOOP
			IF(INPUT(COUNT) = '1') THEN
				tempSUM := tempSUM + 1;
			END IF;
		END LOOP;
			
		SUM <= (2 * tempSUM) - N;
		DONE <= '1';

	END PROCESS;

END RTL;