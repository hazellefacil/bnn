library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity address_counter is
  port(
  
		);
end address_counter;

-- Architecture part of the description

architecture behavioural of address_counter is


begin
	
end behavioural;