library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity part of the description.  Describes inputs and outputs

entity prevariance is
  port(
  
		);
end prevariance;

-- Architecture part of the description

architecture behavioural of prevariance is


begin
	
end behavioural;